//

module demux_32_8(
	input [31:0]		din,
	input [7:0]			selector,
	output reg [7:0]	dout
);
	
	
	always @(*)
		begin
			case((din))
				
				
			endcase
		
		end